module HexHELO( input [0:2] C, output [0:6] Hex);

//Should assign HELO to 0,1,2,3 respectively
assign Hex[0]=  (~C[0]&~C[1]&~C[2])|
			     //( C[0]&~C[1]&~C[2])|
			       (~C[0]& C[1]&~C[2])|
			     //( C[0]& C[1]&~C[2])|
			       (~C[0]&~C[1]& C[2])|
			       ( C[0]&~C[1]& C[2])|
			       (~C[0]& C[1]& C[2])|
			       ( C[0]& C[1]& C[2]);
assign Hex[1]=//(~C[0]&~C[1]&~C[2])|
			       ( C[0]&~C[1]&~C[2])|
			       (~C[0]& C[1]&~C[2])|
			     //( C[0]& C[1]&~C[2])|
			       (~C[0]&~C[1]& C[2])|
			       ( C[0]&~C[1]& C[2])|
			       (~C[0]& C[1]& C[2])|
			       ( C[0]& C[1]& C[2]);
assign Hex[2]=// (~C[0]&~C[1]&~C[2])|
			       ( C[0]&~C[1]&~C[2])|
			       (~C[0]& C[1]&~C[2])|
			     //( C[0]& C[1]&~C[2])|
			       (~C[0]&~C[1]& C[2])|
			       ( C[0]&~C[1]& C[2])|
			       (~C[0]& C[1]& C[2])|
			       ( C[0]& C[1]& C[2]);
assign Hex[3]=  (~C[0]&~C[1]&~C[2])|
			     //( C[0]&~C[1]&~C[2])|
			     //(~C[0]& C[1]&~C[2])|
			     //( C[0]& C[1]&~C[2])|
			       (~C[0]&~C[1]& C[2])|
			       ( C[0]&~C[1]& C[2])|
			       (~C[0]& C[1]& C[2])|
			       ( C[0]& C[1]& C[2]);
assign Hex[4]=//(~C[0]&~C[1]&~C[2])|
			     //( C[0]&~C[1]&~C[2])|
			     //(~C[0]& C[1]&~C[2])|
			     //( C[0]& C[1]&~C[2])|
			       (~C[0]&~C[1]& C[2])|
			       ( C[0]&~C[1]& C[2])|
			       (~C[0]& C[1]& C[2])|
			       ( C[0]& C[1]& C[2]);
assign Hex[5]=//(~C[0]&~C[1]&~C[2])|
			     //( C[0]&~C[1]&~C[2])|
			     //(~C[0]& C[1]&~C[2])|
			     //( C[0]& C[1]&~C[2])|
			       (~C[0]&~C[1]& C[2])|
			       ( C[0]&~C[1]& C[2])|
			       (~C[0]& C[1]& C[2])|
			       ( C[0]& C[1]& C[2]);
assign Hex[6]=//(~C[0]&~C[1]&~C[2])|
			     //( C[0]&~C[1]&~C[2])|
			       (~C[0]& C[1]&~C[2])|
			       ( C[0]& C[1]&~C[2])|
			       (~C[0]&~C[1]& C[2])|
			       ( C[0]&~C[1]& C[2])|
			       (~C[0]& C[1]& C[2])|
			       ( C[0]& C[1]& C[2]);


endmodule
