//Written by:Spencer Sawyer


module HexHEXd( input [3:0] C, output [0:6] Hex);

//Should assign HELO to 0,1,2,3 respectively
assign Hex[0]=//(~C[0]&~C[1]&~C[2])&~C[3]| //0
			       ( C[0]&~C[1]&~C[2])&~C[3]| //1
			     //(~C[0]& C[1]&~C[2])&~C[3]| //2
			     //( C[0]& C[1]&~C[2])&~C[3]| //3
			       (~C[0]&~C[1]& C[2])&~C[3]| //4
			     //( C[0]&~C[1]& C[2])&~C[3]| //5
//			       (~C[0]& C[1]& C[2])&~C[3]| //6
//			       ( C[0]& C[1]& C[2])&~C[3]| //7
//					 (~C[0]&~C[1]&~C[2])& C[3]| //8
//			       ( C[0]&~C[1]&~C[2])& C[3]| //9
//			       (~C[0]& C[1]&~C[2])& C[3]| //A
			       ( C[0]& C[1]&~C[2])& C[3]| //B
//			       (~C[0]&~C[1]& C[2])& C[3]| //C
			       ( C[0]&~C[1]& C[2])& C[3]; //D
//			       (~C[0]& C[1]& C[2])& C[3]| //E
//			       ( C[0]& C[1]& C[2])& C[3]; //F
					 
					 
					 
assign Hex[1]=//(~C[0]&~C[1]&~C[2])&~C[3]| //0
			     //( C[0]&~C[1]&~C[2])&~C[3]| //1
			     //(~C[0]& C[1]&~C[2])&~C[3]| //2
			     //( C[0]& C[1]&~C[2])&~C[3]| //3
			     //(~C[0]&~C[1]& C[2])&~C[3]| //4
			       ( C[0]&~C[1]& C[2])&~C[3]| //5
			       (~C[0]& C[1]& C[2])&~C[3]| //6
//			       ( C[0]& C[1]& C[2])&~C[3]| //7
//					 (~C[0]&~C[1]&~C[2])& C[3]| //8
//			       ( C[0]&~C[1]&~C[2])& C[3]| //9
//			       (~C[0]& C[1]&~C[2])& C[3]| //A
			       ( C[0]& C[1]&~C[2])& C[3]| //B
			       (~C[0]&~C[1]& C[2])& C[3]| //C
//			       ( C[0]&~C[1]& C[2])& C[3]| //D
			       (~C[0]& C[1]& C[2])& C[3]| //E
			       ( C[0]& C[1]& C[2])& C[3]; //F
					 
					 
					 
assign Hex[2]=//(~C[0]&~C[1]&~C[2])&~C[3]| //0
			     //( C[0]&~C[1]&~C[2])&~C[3]| //1
			       (~C[0]& C[1]&~C[2])&~C[3]| //2
			     //( C[0]& C[1]&~C[2])&~C[3]| //3
			     //(~C[0]&~C[1]& C[2])&~C[3]| //4
			     //( C[0]&~C[1]& C[2])&~C[3]| //5
//			       (~C[0]& C[1]& C[2])&~C[3]| //6
//			       ( C[0]& C[1]& C[2])&~C[3]| //7
//					 (~C[0]&~C[1]&~C[2])& C[3]| //8
//			       ( C[0]&~C[1]&~C[2])& C[3]| //9
//			       (~C[0]& C[1]&~C[2])& C[3]| //A
//			       ( C[0]& C[1]&~C[2])& C[3]| //B
			       (~C[0]&~C[1]& C[2])& C[3]| //C
//			       ( C[0]&~C[1]& C[2])& C[3]| //D
			       (~C[0]& C[1]& C[2])& C[3]| //E
			       ( C[0]& C[1]& C[2])& C[3]; //F
					 
					 
					 
assign Hex[3]=//(~C[0]&~C[1]&~C[2])&~C[3]| //0
			       ( C[0]&~C[1]&~C[2])&~C[3]| //1
			     //(~C[0]& C[1]&~C[2])&~C[3]| //2
			     //( C[0]& C[1]&~C[2])&~C[3]| //3
			       (~C[0]&~C[1]& C[2])&~C[3]| //4
//			       ( C[0]&~C[1]& C[2])&~C[3]| //5
//			       (~C[0]& C[1]& C[2])&~C[3]| //6
			       ( C[0]& C[1]& C[2])&~C[3]| //7
//					 (~C[0]&~C[1]&~C[2])& C[3]| //8
//			       ( C[0]&~C[1]&~C[2])& C[3]| //9
			       (~C[0]& C[1]&~C[2])& C[3]| //A
//			       ( C[0]& C[1]&~C[2])& C[3]| //B
//			       (~C[0]&~C[1]& C[2])& C[3]| //C
//			       ( C[0]&~C[1]& C[2])& C[3]| //D
//			       (~C[0]& C[1]& C[2])& C[3]| //E
			       ( C[0]& C[1]& C[2])& C[3]; //F
					 
					 
					 
assign Hex[4]=//(~C[0]&~C[1]&~C[2])&~C[3]| //0
			       ( C[0]&~C[1]&~C[2])&~C[3]| //1
			     //(~C[0]& C[1]&~C[2])&~C[3]| //2
			       ( C[0]& C[1]&~C[2])&~C[3]| //3
			       (~C[0]&~C[1]& C[2])&~C[3]| //4
			       ( C[0]&~C[1]& C[2])&~C[3]| //5
//			       (~C[0]& C[1]& C[2])&~C[3]| //6
			       ( C[0]& C[1]& C[2])&~C[3]| //7
//					 (~C[0]&~C[1]&~C[2])& C[3]| //8
			       ( C[0]&~C[1]&~C[2])& C[3]; //9
//			       (~C[0]& C[1]&~C[2])& C[3]| //A
//			       ( C[0]& C[1]&~C[2])& C[3]| //B
//			       (~C[0]&~C[1]& C[2])& C[3]| //C
//			       ( C[0]&~C[1]& C[2])& C[3]| //D
//			       (~C[0]& C[1]& C[2])& C[3]| //E
//			       ( C[0]& C[1]& C[2])& C[3]; //F
					 
					 
assign Hex[5]=//(~C[0]&~C[1]&~C[2])&~C[3]| //0
			       ( C[0]&~C[1]&~C[2])&~C[3]| //1
			       (~C[0]& C[1]&~C[2])&~C[3]| //2
			       ( C[0]& C[1]&~C[2])&~C[3]| //3
//			       (~C[0]&~C[1]& C[2])&~C[3]| //4
//			       ( C[0]&~C[1]& C[2])&~C[3]| //5
//			       (~C[0]& C[1]& C[2])&~C[3]| //6
			       ( C[0]& C[1]& C[2])&~C[3]| //7
//					 (~C[0]&~C[1]&~C[2])& C[3]| //8
//			       ( C[0]&~C[1]&~C[2])& C[3]| //9
//			       (~C[0]& C[1]&~C[2])& C[3]| //A
//			       ( C[0]& C[1]&~C[2])& C[3]| //B
//			       (~C[0]&~C[1]& C[2])& C[3]| //C
			       ( C[0]&~C[1]& C[2])& C[3]; //D
//			       (~C[0]& C[1]& C[2])& C[3]| //E
//			       ( C[0]& C[1]& C[2])& C[3]; //F

					 
assign Hex[6]=  (~C[0]&~C[1]&~C[2])&~C[3]| //0
			       ( C[0]&~C[1]&~C[2])&~C[3]| //1
			     //(~C[0]& C[1]&~C[2])&~C[3]| //2
			     //( C[0]& C[1]&~C[2])&~C[3]| //3
			     //(~C[0]&~C[1]& C[2])&~C[3]| //4
//			       ( C[0]&~C[1]& C[2])&~C[3]| //5
//			       (~C[0]& C[1]& C[2])&~C[3]| //6
			       ( C[0]& C[1]& C[2])&~C[3]| //7
//					 (~C[0]&~C[1]&~C[2])& C[3]| //8
//			       ( C[0]&~C[1]&~C[2])& C[3]| //9
//			       (~C[0]& C[1]&~C[2])& C[3]| //A
//			       ( C[0]& C[1]&~C[2])& C[3]| //B
			       (~C[0]&~C[1]& C[2])& C[3]; //C
//			       ( C[0]&~C[1]& C[2])& C[3]| //D
//			       (~C[0]& C[1]& C[2])& C[3]| //E
//			       ( C[0]& C[1]& C[2])& C[3]; //F


endmodule
